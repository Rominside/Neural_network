// -------------------------------------------------------------------
// @author ochir
// @copyright (C) 2023, <COMPANY>
//
// Created : 04. окт. 2023 1:07
//-------------------------------------------------------------------
module Layer ();



endmodule : Layer